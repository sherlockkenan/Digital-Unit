/*module y86decode(y86_inst,mips_inst);
input[63:0] y86_inst;
output[31:0] mips_inst;

//assign mips_inst=y86_inst[63:32];  
always @ (*)
case 
;
endcase
endmodule*/